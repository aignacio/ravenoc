`ifndef _RAVENOC_PKG_
  `define _RAVENOC_PKG_
  package ravenoc_pkg;
    `include  "ravenoc_defines.svh"
    `include  "ravenoc_structs.svh"
    `include  "ravenoc_axi_fnc.svh"
  endpackage
`endif
