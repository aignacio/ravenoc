`ifndef _ravenoc_pkg_
  `define _ravenoc_pkg_
  package ravenoc_pkg;
    //`include  "ravenoc_defines.svh"
    `include  "ravenoc_structs.svh"
  endpackage
`endif
