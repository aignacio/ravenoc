`ifndef _ravenoc_defines_
  `define _ravenoc_defines_
  localparam  FLIT_WIDTH  = 34;  // Flit width in bits
  localparam  N_VIRT_CHN  = 2;   // Number of virtual channels
`endif
